*** SPICE deck for cell 8-Bit-RCA{sch} from library ripple_carry_adders
*** Created on Sat Oct 12, 2019 12:53:54
*** Last revised on Sat Oct 12, 2019 14:53:53
*** Written on Sat Oct 12, 2019 14:53:59 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT ripple_carry_adders__FullAdder FROM CELL FullAdder{sch}
.SUBCKT ripple_carry_adders__FullAdder A B CarryOut Cin Sum
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@29 Cin net@23 gnd NMOS L=0.35U W=0.875U
Mnmos@1 net@23 A gnd gnd NMOS L=0.35U W=0.875U
Mnmos@2 net@23 B gnd gnd NMOS L=0.35U W=0.875U
Mnmos@3 net@29 A net@25 gnd NMOS L=0.35U W=0.875U
Mnmos@4 net@25 B gnd gnd NMOS L=0.35U W=0.875U
Mnmos@5 CarryOut net@29 gnd gnd NMOS L=0.35U W=0.875U
Mnmos@6 net@74 net@29 net@81 gnd NMOS L=0.35U W=0.875U
Mnmos@7 net@81 A gnd gnd NMOS L=0.35U W=0.875U
Mnmos@8 net@81 B gnd gnd NMOS L=0.35U W=0.875U
Mnmos@9 net@81 Cin gnd gnd NMOS L=0.35U W=0.875U
Mnmos@10 net@74 A net@100 gnd NMOS L=0.35U W=0.875U
Mnmos@11 net@100 B net@101 gnd NMOS L=0.35U W=0.875U
Mnmos@12 net@101 Cin gnd gnd NMOS L=0.35U W=0.875U
Mnmos@13 Sum net@74 gnd gnd NMOS L=0.35U W=0.875U
Mpmos@0 vdd A net@0 vdd PMOS L=0.35U W=1.75U
Mpmos@1 net@0 A net@18 vdd PMOS L=0.35U W=1.75U
Mpmos@2 vdd B net@0 vdd PMOS L=0.35U W=1.75U
Mpmos@3 net@0 Cin net@29 vdd PMOS L=0.35U W=1.75U
Mpmos@4 net@18 B net@29 vdd PMOS L=0.35U W=1.75U
Mpmos@5 vdd net@29 CarryOut vdd PMOS L=0.35U W=1.75U
Mpmos@6 net@59 net@29 net@74 vdd PMOS L=0.35U W=1.75U
Mpmos@7 vdd A net@59 vdd PMOS L=0.35U W=1.75U
Mpmos@8 vdd B net@59 vdd PMOS L=0.35U W=1.75U
Mpmos@9 vdd Cin net@59 vdd PMOS L=0.35U W=1.75U
Mpmos@10 net@59 A net@72 vdd PMOS L=0.35U W=1.75U
Mpmos@11 net@72 B net@73 vdd PMOS L=0.35U W=1.75U
Mpmos@12 net@73 Cin net@74 vdd PMOS L=0.35U W=1.75U
Mpmos@13 vdd net@74 Sum vdd PMOS L=0.35U W=1.75U
.ENDS ripple_carry_adders__FullAdder

.global gnd vdd

*** TOP LEVEL CELL: 8-Bit-RCA{sch}
XFullAdde@9 A0 B0 net@41 Cin Sum0 ripple_carry_adders__FullAdder
XFullAdde@10 A1 B1 net@47 net@41 Sum1 ripple_carry_adders__FullAdder
XFullAdde@11 A2 B2 net@52 net@47 Sum2 ripple_carry_adders__FullAdder
XFullAdde@12 A3 B3 net@58 net@52 Sum3 ripple_carry_adders__FullAdder
XFullAdde@13 A4 B4 net@62 net@58 Sum4 ripple_carry_adders__FullAdder
XFullAdde@14 A5 B5 net@67 net@62 Sum5 ripple_carry_adders__FullAdder
XFullAdde@15 A6 B6 net@72 net@67 Sum6 ripple_carry_adders__FullAdder
XFullAdde@16 A7 B7 Cout net@72 Sum7 ripple_carry_adders__FullAdder

* Spice Code nodes in cell cell '8-Bit-RCA{sch}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
Vin A0 0 DC 0
Vin2 A1 0 DC 0
Vin3 A2 0 DC 3.3
Vin4 A3 0 DC 3.3
Vin5 A4 0 DC 0
Vin6 A5 0 DC 0
Vin7 A6 0 DC 0
Vin8 A7 0 DC 0
Vin9 B0 0 DC 3.3
Vin10 B1 0 DC 0
Vin11 B2 0 DC 3.3
Vin12 B3 0 DC 3.3
Vin13 B4 0 DC 0
Vin14 B5 0 DC 0
Vin15 B6 0 DC 0
Vin16 B7 0 DC 0
Vin17 Cin 0 DC 0
.TRAN 0 100n
.include C:\Users\kille\Desktop\Electric\C5_models.txt
.END
