*** SPICE deck for cell xyzw{sch} from library Homework_4
*** Created on Sat Nov 02, 2019 20:31:47
*** Last revised on Sat Nov 02, 2019 23:01:06
*** Written on Sat Nov 02, 2019 23:06:15 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: Homework_4:xyzw{sch}
Ccap@0 gnd net@14 5p
Mnmos@0 net@9 Clock gnd gnd NMOS L=0.35U W=0.875U
Mnmos@2 net@14 X net@2 gnd NMOS L=0.35U W=0.875U
Mnmos@3 net@2 Y net@9 gnd NMOS L=0.35U W=0.875U
Mnmos@4 net@14 X net@6 gnd NMOS L=0.35U W=0.875U
Mnmos@5 net@6 Z net@9 gnd NMOS L=0.35U W=0.875U
Mnmos@6 net@6 W net@9 gnd NMOS L=0.35U W=0.875U
Mpmos@0 vdd Clock net@14 vdd PMOS L=0.35U W=1.75U

* Spice Code nodes in cell cell 'Homework_4:xyzw{sch}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
Vin X 0 dc 3.3
Vin1 Z 0 dc 3.3
Vin2 W 0 dc 3.3
Vin3 Y 0 dc PULSE (0 1 0 0.1n 0.1n 0.5s 1s)
Vin4 Clock 0 dc PULSE (0 1 0 0.1n 0.1n 1s 2s)
cload F out 0 5pF
.TRAN 0 6s
.include C:\Users\kille\Desktop\Electric\C5_models.txt
.END
